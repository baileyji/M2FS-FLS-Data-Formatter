------------------------------------------------------------
-- VHDL M2FS_FLS_Data_Formatter_FPGA_8_14_2012
-- 2012 10 19 13 56 2
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2004 Altium Limited"
------------------------------------------------------------

------------------------------------------------------------
-- VHDL M2FS_FLS_Data_Formatter_FPGA_8_14_2012
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity M2FS_FLS_Data_Formatter_FPGA_8_14_2012 Is
  attribute MacroCell : boolean;

End M2FS_FLS_Data_Formatter_FPGA_8_14_2012;
------------------------------------------------------------

------------------------------------------------------------
architecture structure of M2FS_FLS_Data_Formatter_FPGA_8_14_2012 is


begin
end structure;
------------------------------------------------------------

